module BIOS
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=10)
(
	input [(ADDR_WIDTH-1):0] addr,
	input clk, 
	output reg [(DATA_WIDTH-1):0] q
);
	reg [DATA_WIDTH-1:0] BIOS[2**ADDR_WIDTH-1:0];

	initial
	begin: INIT
BIOS[0] = 32'b01101_11101_00000_00000000000000000;
BIOS[1] = 32'b10101_000000000000000000000000010;
BIOS[2] = 32'b01101_00001_00000_00000000001100011;
BIOS[3] = 32'b00000_10010_00001_00000_000000000000;
BIOS[4] = 32'b01100_10010_00000_00000_000000000000;
BIOS[5] = 32'b01101_00011_00000_00000000001100010;
BIOS[6] = 32'b00000_10010_00011_00000_000000000000;
BIOS[7] = 32'b01100_10010_00000_00000_000000000000;
BIOS[8] = 32'b01101_00101_00000_00000000000000001;
BIOS[9] = 32'b00000_10010_00101_00000_000000000000;
BIOS[10] = 32'b01101_00110_00000_00000000000000000;
BIOS[11] = 32'b00000_10011_00110_00000_000000000000;
BIOS[12] = 32'b01101_00111_00000_00000000000011000;
BIOS[13] = 32'b00000_10100_00111_00000_000000000000;
BIOS[14] = 32'b11111_10010_10011_10100_000000000000;
BIOS[15] = 32'b01101_01001_00000_00000000000010001;
BIOS[16] = 32'b00000_10010_01001_00000_000000000000;
BIOS[17] = 32'b01101_01010_00000_00000000000000000;
BIOS[18] = 32'b00000_10011_01010_00000_000000000000;
BIOS[19] = 32'b01101_01011_00000_00000000000011000;
BIOS[20] = 32'b00000_10100_01011_00000_000000000000;
BIOS[21] = 32'b11110_10010_10011_10100_000000000000;
BIOS[22] = 32'b01100_00001_00000_00000_000000000000;
BIOS[23] = 32'b11001_000000000000000000000000000;
	end

	always @ (posedge clk)
	begin
		q <= BIOS[addr];
	end

endmodule
